module keySchedule(
    );


endmodule
