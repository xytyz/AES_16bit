module LUT_verilog( 
	output reg [7:0]outp, 
	input [7:0] inp
    );
	
	always @(inp) begin
		case(inp)
			8'h00: outp<= 8'h63;
			8'h01: outp<= 8'h7c;
			8'h02: outp<= 8'h77;
			8'h03: outp<= 8'h7b;
			8'h04: outp<= 8'hf2;
			8'h05: outp<= 8'h6b;
			8'h06: outp<= 8'h6f;
			8'h07: outp<= 8'hc5;
			8'h08: outp<= 8'h30;
			8'h09: outp<= 8'h01;
			8'h0a: outp<= 8'h67;
			8'h0b: outp<= 8'h2b;
			8'h0c: outp<= 8'hfe;
			8'h0d: outp<= 8'hd7;
			8'h0e: outp<= 8'hab;
			8'h0f: outp<= 8'h76;
			8'h10: outp<= 8'hca;
			8'h11: outp<= 8'h82;
			8'h12: outp<= 8'hc9;
			8'h13: outp<= 8'h7d;
			8'h14: outp<= 8'hfa;
			8'h15: outp<= 8'h59;
			8'h16: outp<= 8'h47;
			8'h17: outp<= 8'hf0;
			8'h18: outp<= 8'had;
			8'h19: outp<= 8'hd4;
			8'h1a: outp<= 8'ha2;
			8'h1b: outp<= 8'haf;
			8'h1c: outp<= 8'h9c;
			8'h1d: outp<= 8'ha4;
			8'h1e: outp<= 8'h72;
			8'h1f: outp<= 8'hc0;
			8'h20: outp<= 8'hb7;
			8'h21: outp<= 8'hfd;
			8'h22: outp<= 8'h93;
			8'h23: outp<= 8'h26;
			8'h24: outp<= 8'h36;
			8'h25: outp<= 8'h3f;
			8'h26: outp<= 8'hf7;
			8'h27: outp<= 8'hcc;
			8'h28: outp<= 8'h34;
			8'h29: outp<= 8'ha5;
			8'h2a: outp<= 8'he5;
			8'h2b: outp<= 8'hf1;
			8'h2c: outp<= 8'h71;
			8'h2d: outp<= 8'hd8;
			8'h2e: outp<= 8'h31;
			8'h2f: outp<= 8'h15;
			8'h30: outp<= 8'h04;
			8'h31: outp<= 8'hc7;
			8'h32: outp<= 8'h23;
			8'h33: outp<= 8'hc3;
			8'h34: outp<= 8'h18;
			8'h35: outp<= 8'h96;
			8'h36: outp<= 8'h05;
			8'h37: outp<= 8'h9a;
			8'h38: outp<= 8'h07;
			8'h39: outp<= 8'h12;
			8'h3a: outp<= 8'h80;
			8'h3b: outp<= 8'he2;
			8'h3c: outp<= 8'heb;
			8'h3d: outp<= 8'h27;
			8'h3e: outp<= 8'hb2;
			8'h3f: outp<= 8'h75;
			8'h40: outp<= 8'h09;
			8'h41: outp<= 8'h83;
			8'h42: outp<= 8'h2c;
			8'h43: outp<= 8'h1a;
			8'h44: outp<= 8'h1b;
			8'h45: outp<= 8'h6e;
			8'h46: outp<= 8'h5a;
			8'h47: outp<= 8'ha0;
			8'h48: outp<= 8'h52;
			8'h49: outp<= 8'h3b;
			8'h4a: outp<= 8'hd6;
			8'h4b: outp<= 8'hb3;
			8'h4c: outp<= 8'h29;
			8'h4d: outp<= 8'he3;
			8'h4e: outp<= 8'h2f;
			8'h4f: outp<= 8'h84;
			8'h50: outp<= 8'h53;
			8'h51: outp<= 8'hd1;
			8'h52: outp<= 8'h00;
			8'h53: outp<= 8'hed;
			8'h54: outp<= 8'h20;
			8'h55: outp<= 8'hfc;
			8'h56: outp<= 8'hb1;
			8'h57: outp<= 8'h5b;
			8'h58: outp<= 8'h6a;
			8'h59: outp<= 8'hcb;
			8'h5a: outp<= 8'hbe;
			8'h5b: outp<= 8'h39;
			8'h5c: outp<= 8'h4a;
			8'h5d: outp<= 8'h4c;
			8'h5e: outp<= 8'h58;
			8'h5f: outp<= 8'hcf;
			8'h60: outp<= 8'hd0;
			8'h61: outp<= 8'hef;
			8'h62: outp<= 8'haa;
			8'h63: outp<= 8'hfb;
			8'h64: outp<= 8'h43;
			8'h65: outp<= 8'h4d;
			8'h66: outp<= 8'h33;
			8'h67: outp<= 8'h85;
			8'h68: outp<= 8'h45;
			8'h69: outp<= 8'hf9;
			8'h6a: outp<= 8'h02;
			8'h6b: outp<= 8'h7f;
			8'h6c: outp<= 8'h50;
			8'h6d: outp<= 8'h3c;
			8'h6e: outp<= 8'h9f;
			8'h6f: outp<= 8'ha8;
			8'h70: outp<= 8'h51;
			8'h71: outp<= 8'ha3;
			8'h72: outp<= 8'h40;
			8'h73: outp<= 8'h8f;
			8'h74: outp<= 8'h92;
			8'h75: outp<= 8'h9d;
			8'h76: outp<= 8'h38;
			8'h77: outp<= 8'hf5;
			8'h78: outp<= 8'hbc;
			8'h79: outp<= 8'hb6;
			8'h7a: outp<= 8'hda;
			8'h7b: outp<= 8'h21;
			8'h7c: outp<= 8'h10;
			8'h7d: outp<= 8'hff;
			8'h7e: outp<= 8'hf3;
			8'h7f: outp<= 8'hd2;
			8'h80: outp<= 8'hcd;
			8'h81: outp<= 8'h0c;
			8'h82: outp<= 8'h13;
			8'h83: outp<= 8'hec;
			8'h84: outp<= 8'h5f;
			8'h85: outp<= 8'h97;
			8'h86: outp<= 8'h44;
			8'h87: outp<= 8'h17;
			8'h88: outp<= 8'hc4;
			8'h89: outp<= 8'ha7;
			8'h8a: outp<= 8'h7e;
			8'h8b: outp<= 8'h3d;
			8'h8c: outp<= 8'h64;
			8'h8d: outp<= 8'h5d;
			8'h8e: outp<= 8'h19;
			8'h8f: outp<= 8'h73;
			8'h90: outp<= 8'h60;
			8'h91: outp<= 8'h81;
			8'h92: outp<= 8'h4f;
			8'h93: outp<= 8'hdc;
			8'h94: outp<= 8'h22;
			8'h95: outp<= 8'h2a;
			8'h96: outp<= 8'h90;
			8'h97: outp<= 8'h88;
			8'h98: outp<= 8'h46;
			8'h99: outp<= 8'hee;
			8'h9a: outp<= 8'hb8;
			8'h9b: outp<= 8'h14;
			8'h9c: outp<= 8'hde;
			8'h9d: outp<= 8'h5e;
			8'h9e: outp<= 8'h0b;
			8'h9f: outp<= 8'hdb;
			8'ha0: outp<= 8'he0;
			8'ha1: outp<= 8'h32;
			8'ha2: outp<= 8'h3a;
			8'ha3: outp<= 8'h0a;
			8'ha4: outp<= 8'h49;
			8'ha5: outp<= 8'h06;
			8'ha6: outp<= 8'h24;
			8'ha7: outp<= 8'h5c;
			8'ha8: outp<= 8'hc2;
			8'ha9: outp<= 8'hd3;
			8'haa: outp<= 8'hac;
			8'hab: outp<= 8'h62;
			8'hac: outp<= 8'h91;
			8'had: outp<= 8'h95;
			8'hae: outp<= 8'he4;
			8'haf: outp<= 8'h79;
			8'hb0: outp<= 8'he7;
			8'hb1: outp<= 8'hc8;
			8'hb2: outp<= 8'h37;
			8'hb3: outp<= 8'h6d;
			8'hb4: outp<= 8'h8d;
			8'hb5: outp<= 8'hd5;
			8'hb6: outp<= 8'h4e;
			8'hb7: outp<= 8'ha9;
			8'hb8: outp<= 8'h6c;
			8'hb9: outp<= 8'h56;
			8'hba: outp<= 8'hf4;
			8'hbb: outp<= 8'hea;
			8'hbc: outp<= 8'h65;
			8'hbd: outp<= 8'h7a;
			8'hbe: outp<= 8'hae;
			8'hbf: outp<= 8'h08;
			8'hc0: outp<= 8'hba;
			8'hc1: outp<= 8'h78;
			8'hc2: outp<= 8'h25;
			8'hc3: outp<= 8'h2e;
			8'hc4: outp<= 8'h1c;
			8'hc5: outp<= 8'ha6;
			8'hc6: outp<= 8'hb4;
			8'hc7: outp<= 8'hc6;
			8'hc8: outp<= 8'he8;
			8'hc9: outp<= 8'hdd;
			8'hca: outp<= 8'h74;
			8'hcb: outp<= 8'h1f;
			8'hcc: outp<= 8'h4b;
			8'hcd: outp<= 8'hbd;
			8'hce: outp<= 8'h8b;
			8'hcf: outp<= 8'h8a;
			8'hd0: outp<= 8'h70;
			8'hd1: outp<= 8'h3e;
			8'hd2: outp<= 8'hb5;
			8'hd3: outp<= 8'h66;
			8'hd4: outp<= 8'h48;
			8'hd5: outp<= 8'h03;
			8'hd6: outp<= 8'hf6;
			8'hd7: outp<= 8'h0e;
			8'hd8: outp<= 8'h61;
			8'hd9: outp<= 8'h35;
			8'hda: outp<= 8'h57;
			8'hdb: outp<= 8'hb9;
			8'hdc: outp<= 8'h86;
			8'hdd: outp<= 8'hc1;
			8'hde: outp<= 8'h1d;
			8'hdf: outp<= 8'h9e;
			8'he0: outp<= 8'he1;
			8'he1: outp<= 8'hf8;
			8'he2: outp<= 8'h98;
			8'he3: outp<= 8'h11;
			8'he4: outp<= 8'h69;
			8'he5: outp<= 8'hd9;
			8'he6: outp<= 8'h8e;
			8'he7: outp<= 8'h94;
			8'he8: outp<= 8'h9b;
			8'he9: outp<= 8'h1e;
			8'hea: outp<= 8'h87;
			8'heb: outp<= 8'he9;
			8'hec: outp<= 8'hce;
			8'hed: outp<= 8'h55;
			8'hee: outp<= 8'h28;
			8'hef: outp<= 8'hdf;
			8'hf0: outp<= 8'h8c;
			8'hf1: outp<= 8'ha1;
			8'hf2: outp<= 8'h89;
			8'hf3: outp<= 8'h0d;
			8'hf4: outp<= 8'hbf;
			8'hf5: outp<= 8'he6;
			8'hf6: outp<= 8'h42;
			8'hf7: outp<= 8'h68;
			8'hf8: outp<= 8'h41;
			8'hf9: outp<= 8'h99;
			8'hfa: outp<= 8'h2d;
			8'hfb: outp<= 8'h0f;
			8'hfc: outp<= 8'hb0;
			8'hfd: outp<= 8'h54;
			8'hfe: outp<= 8'hbb;
			8'hff: outp<= 8'h16;
		endcase
	end

endmodule
