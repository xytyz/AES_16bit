module mixCol(
	input [15:0] code,
	output [15:0] altered
    );
	 
assign altered[15]= code[15:0];


endmodule
