module inv_LUT(output reg [7:0] code, input [7:0] inp
    );
	
	always @(inp) begin
		case(inp)
			8'h00: code<= 8'h52;
			8'h01: code<= 8'h09;
			8'h02: code<= 8'h6a;
			8'h03: code<= 8'hd5;
			8'h04: code<= 8'h30;
			8'h05: code<= 8'h36;
			8'h06: code<= 8'ha5;
			8'h07: code<= 8'h38;
			8'h08: code<= 8'hbf;
			8'h09: code<= 8'h40;
			8'h0a: code<= 8'ha3;
			8'h0b: code<= 8'h9e;
			8'h0c: code<= 8'h81;
			8'h0d: code<= 8'hf3;
			8'h0e: code<= 8'hd7;
			8'h0f: code<= 8'hfb;
			8'h10: code<= 8'h7c;
			8'h11: code<= 8'he3;
			8'h12: code<= 8'h39;
			8'h13: code<= 8'h82;
			8'h14: code<= 8'h9b;
			8'h15: code<= 8'h2f;
			8'h16: code<= 8'hff;
			8'h17: code<= 8'h87;
			8'h18: code<= 8'h34;
			8'h19: code<= 8'h8e;
			8'h1a: code<= 8'h43;
			8'h1b: code<= 8'h44;
			8'h1c: code<= 8'hc4;
			8'h1d: code<= 8'hde;
			8'h1e: code<= 8'he9;
			8'h1f: code<= 8'hcb;
			8'h20: code<= 8'h54;
			8'h21: code<= 8'h7b;
			8'h22: code<= 8'h94;
			8'h23: code<= 8'h32;
			8'h24: code<= 8'ha6;
			8'h25: code<= 8'hc2;
			8'h26: code<= 8'h23;
			8'h27: code<= 8'h3d;
			8'h28: code<= 8'hee;
			8'h29: code<= 8'h4c;
			8'h2a: code<= 8'h95;
			8'h2b: code<= 8'h0b;
			8'h2c: code<= 8'h42;
			8'h2d: code<= 8'hfa;
			8'h2e: code<= 8'hc3;
			8'h2f: code<= 8'h4e;
			8'h30: code<= 8'h08;
			8'h31: code<= 8'h2e;
			8'h32: code<= 8'ha1;
			8'h33: code<= 8'h66;
			8'h34: code<= 8'h28;
			8'h35: code<= 8'hd9;
			8'h36: code<= 8'h24;
			8'h37: code<= 8'hb2;
			8'h38: code<= 8'h76;
			8'h39: code<= 8'h5b;
			8'h3a: code<= 8'ha2;
			8'h3b: code<= 8'h49;
			8'h3c: code<= 8'h6d;
			8'h3d: code<= 8'h8b;
			8'h3e: code<= 8'hd1;
			8'h3f: code<= 8'h25;
			8'h40: code<= 8'h72;
			8'h41: code<= 8'hf8;
			8'h42: code<= 8'hf6;
			8'h43: code<= 8'h64;
			8'h44: code<= 8'h86;
			8'h45: code<= 8'h68;
			8'h46: code<= 8'h98;
			8'h47: code<= 8'h16;
			8'h48: code<= 8'hd4;
			8'h49: code<= 8'ha4;
			8'h4a: code<= 8'h5c;
			8'h4b: code<= 8'hcc;
			8'h4c: code<= 8'h5d;
			8'h4d: code<= 8'h65;
			8'h4e: code<= 8'hb6;
			8'h4f: code<= 8'h92;
			8'h50: code<= 8'h6c;
			8'h51: code<= 8'h70;
			8'h52: code<= 8'h48;
			8'h53: code<= 8'h50;
			8'h54: code<= 8'hfd;
			8'h55: code<= 8'hed;
			8'h56: code<= 8'hb9;
			8'h57: code<= 8'hda;
			8'h58: code<= 8'h5e;
			8'h59: code<= 8'h15;
			8'h5a: code<= 8'h46;
			8'h5b: code<= 8'h57;
			8'h5c: code<= 8'ha7;
			8'h5d: code<= 8'h8d;
			8'h5e: code<= 8'h9d;
			8'h5f: code<= 8'h84;
			8'h60: code<= 8'h90;
			8'h61: code<= 8'hd8;
			8'h62: code<= 8'hab;
			8'h63: code<= 8'h00;
			8'h64: code<= 8'h8c;
			8'h65: code<= 8'hbc;
			8'h66: code<= 8'hd3;
			8'h67: code<= 8'h0a;
			8'h68: code<= 8'hf7;
			8'h69: code<= 8'he4;
			8'h6a: code<= 8'h58;
			8'h6b: code<= 8'h05;
			8'h6c: code<= 8'hb8;
			8'h6d: code<= 8'hb3;
			8'h6e: code<= 8'h45;
			8'h6f: code<= 8'h06;
			8'h70: code<= 8'hd0;
			8'h71: code<= 8'h2c;
			8'h72: code<= 8'h1e;
			8'h73: code<= 8'h8f;
			8'h74: code<= 8'hca;
			8'h75: code<= 8'h3f;
			8'h76: code<= 8'h0f;
			8'h77: code<= 8'h02;
			8'h78: code<= 8'hc1;
			8'h79: code<= 8'haf;
			8'h7a: code<= 8'hbd;
			8'h7b: code<= 8'h03;
			8'h7c: code<= 8'h01;
			8'h7d: code<= 8'h13;
			8'h7e: code<= 8'h8a;
			8'h7f: code<= 8'h6b;
			8'h80: code<= 8'h3a;
			8'h81: code<= 8'h91;
			8'h82: code<= 8'h11;
			8'h83: code<= 8'h41;
			8'h84: code<= 8'h4f;
			8'h85: code<= 8'h67;
			8'h86: code<= 8'hdc;
			8'h87: code<= 8'hea;
			8'h88: code<= 8'h97;
			8'h89: code<= 8'hf2;
			8'h8a: code<= 8'hcf;
			8'h8b: code<= 8'hce;
			8'h8c: code<= 8'hf0;
			8'h8d: code<= 8'hb4;
			8'h8e: code<= 8'he6;
			8'h8f: code<= 8'h73;
			8'h90: code<= 8'h96;
			8'h91: code<= 8'hac;
			8'h92: code<= 8'h74;
			8'h93: code<= 8'h22;
			8'h94: code<= 8'he7;
			8'h95: code<= 8'had;
			8'h96: code<= 8'h35;
			8'h97: code<= 8'h85;
			8'h98: code<= 8'he2;
			8'h99: code<= 8'hf9;
			8'h9a: code<= 8'h37;
			8'h9b: code<= 8'he8;
			8'h9c: code<= 8'h1c;
			8'h9d: code<= 8'h75;
			8'h9e: code<= 8'hdf;
			8'h9f: code<= 8'h6e;
			8'ha0: code<= 8'h47;
			8'ha1: code<= 8'hf1;
			8'ha2: code<= 8'h1a;
			8'ha3: code<= 8'h71;
			8'ha4: code<= 8'h1d;
			8'ha5: code<= 8'h29;
			8'ha6: code<= 8'hc5;
			8'ha7: code<= 8'h89;
			8'ha8: code<= 8'h6f;
			8'ha9: code<= 8'hb7;
			8'haa: code<= 8'h62;
			8'hab: code<= 8'h0e;
			8'hac: code<= 8'haa;
			8'had: code<= 8'h18;
			8'hae: code<= 8'hbe;
			8'haf: code<= 8'h1b;
			8'hb0: code<= 8'hfc;
			8'hb1: code<= 8'h56;
			8'hb2: code<= 8'h3e;
			8'hb3: code<= 8'h4b;
			8'hb4: code<= 8'hc6;
			8'hb5: code<= 8'hd2;
			8'hb6: code<= 8'h79;
			8'hb7: code<= 8'h20;
			8'hb8: code<= 8'h9a;
			8'hb9: code<= 8'hdb;
			8'hba: code<= 8'hc0;
			8'hbb: code<= 8'hfe;
			8'hbc: code<= 8'h78;
			8'hbd: code<= 8'hcd;
			8'hbe: code<= 8'h5a;
			8'hbf: code<= 8'hf4;
			8'hc0: code<= 8'h1f;
			8'hc1: code<= 8'hdd;
			8'hc2: code<= 8'ha8;
			8'hc3: code<= 8'h33;
			8'hc4: code<= 8'h88;
			8'hc5: code<= 8'h07;
			8'hc6: code<= 8'hc7;
			8'hc7: code<= 8'h31;
			8'hc8: code<= 8'hb1;
			8'hc9: code<= 8'h12;
			8'hca: code<= 8'h10;
			8'hcb: code<= 8'h59;
			8'hcc: code<= 8'h27;
			8'hcd: code<= 8'h80;
			8'hce: code<= 8'hec;
			8'hcf: code<= 8'h5f;
			8'hd0: code<= 8'h60;
			8'hd1: code<= 8'h51;
			8'hd2: code<= 8'h7f;
			8'hd3: code<= 8'ha9;
			8'hd4: code<= 8'h19;
			8'hd5: code<= 8'hb5;
			8'hd6: code<= 8'h4a;
			8'hd7: code<= 8'h0d;
			8'hd8: code<= 8'h2d;
			8'hd9: code<= 8'he5;
			8'hda: code<= 8'h7a;
			8'hdb: code<= 8'h9f;
			8'hdc: code<= 8'h93;
			8'hdd: code<= 8'hc9;
			8'hde: code<= 8'h9c;
			8'hdf: code<= 8'hef;
			8'he0: code<= 8'ha0;
			8'he1: code<= 8'he0;
			8'he2: code<= 8'h3b;
			8'he3: code<= 8'h4d;
			8'he4: code<= 8'hae;
			8'he5: code<= 8'h2a;
			8'he6: code<= 8'hf5;
			8'he7: code<= 8'hb0;
			8'he8: code<= 8'hc8;
			8'he9: code<= 8'heb;
			8'hea: code<= 8'hbb;
			8'heb: code<= 8'h3c;
			8'hec: code<= 8'h83;
			8'hed: code<= 8'h53;
			8'hee: code<= 8'h99;
			8'hef: code<= 8'h61;
			8'hf0: code<= 8'h17;
			8'hf1: code<= 8'h2b;
			8'hf2: code<= 8'h04;
			8'hf3: code<= 8'h7e;
			8'hf4: code<= 8'hba;
			8'hf5: code<= 8'h77;
			8'hf6: code<= 8'hd6;
			8'hf7: code<= 8'h26;
			8'hf8: code<= 8'he1;
			8'hf9: code<= 8'h69;
			8'hfa: code<= 8'h14;
			8'hfb: code<= 8'h63;
			8'hfc: code<= 8'h55;
			8'hfd: code<= 8'h21;
			8'hfe: code<= 8'h0c;
			8'hff: code<= 8'h7d;
			default: code<= 8'h00;
		endcase
	end
endmodule
